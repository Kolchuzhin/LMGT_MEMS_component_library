package initial_160 is

constant mm_1:real:=  0.306735124580E-07;
constant km_1:real:=  23.67780511942;		-- ddE/dq1/dq1 at q1=0.0
constant dm_1:real:=  2.840743666170e-05;	-- Q=30

constant mm_2:real:=  0.201756803926E-07;
constant km_2:real:=  212.6896178680;		-- ddE/dq2/dq2 at q2=0.0
constant dm_2:real:=  6.905036631344e-05;	-- Q=30

constant fi1_1:real:=   1.00000000000    ;
constant fi1_2:real:=   1.00000000000    ;
constant fi2_1:real:=  0.999999560836    ;
constant fi2_2:real:=  0.999998225220    ;

end;
