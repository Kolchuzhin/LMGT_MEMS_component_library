package s_dat_160 is

constant s_type160:integer:=1;
constant s_inve160:integer:=1;
signal s_ord160:real_vector(1 to 3):=( 4.0, 4.0, 0.0 );
signal s_fak160:real_vector(1 to 4):=( 0.114386722375, 0.795085352965, 0.0, 2107.233904 );
constant s_anz160:integer:=      25;
signal s_data160:real_vector(1 to 25):=
(
  0.832702752873E-07,
 -0.140453798427E-14,
  0.429309184785    ,
  0.109391250030E-14,
  0.291985344904    ,
  0.207339774625E-14,
 -0.186971620812E-05,
 -0.152582657928E-13,
  0.124224281759    ,
  0.148706670364E-13,
  0.798129483956E-01,
  0.206229910840E-13,
  0.627255053996E-01,
 -0.205185875145E-13,
  0.153987606242E-05,
 -0.247538941670E-14,
  0.104493898549E-01,
  0.183901764210E-13,
  0.516669367876E-06,
 -0.179097341258E-13,
  0.149282741683E-02,
 -0.189532739990E-13,
  0.143077040992E-06,
  0.189540164009E-13,
  0.216911589898E-08
);

end;
