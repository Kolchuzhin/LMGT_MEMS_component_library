package ca12_dat_160 is

constant ca12_type160:integer:=1;
constant ca12_inve160:integer:=2;
signal ca12_ord160:real_vector(1 to 3):=( 4.0, 4.0, 0.0 );
signal ca12_fak160:real_vector(1 to 4):=( 0.114386722375, 0.795085352965, 0.0, 0.225083783539 );
constant ca12_anz160:integer:=      25;
signal ca12_data160:real_vector(1 to 25):=
(
  0.924864850772    ,
  0.750140219005E-01,
 -0.661841035530E-02,
  0.109715066982E-02,
 -0.215094781164E-03,
 -0.533643405991E-02,
 -0.864001014363E-03,
  0.315112801689E-03,
 -0.103808114827E-03,
  0.301052576502E-04,
 -0.142570841390E-03,
  0.546854159479E-04,
 -0.209086737993E-04,
  0.897245384403E-05,
 -0.318291521927E-05,
  0.160290107930E-05,
 -0.173411215981E-05,
  0.101851559925E-05,
 -0.625232626794E-06,
  0.277844130785E-06,
 -0.774100642402E-07,
  0.824389854108E-07,
 -0.539399052887E-07,
  0.362089073215E-07,
 -0.191260647195E-07
);

end;
