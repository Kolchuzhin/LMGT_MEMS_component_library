-- Analytical based model of a micro-mirror
-- coming soon ...
