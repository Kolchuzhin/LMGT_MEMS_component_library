-- Analytical based model of a micro-electro-mechanical transducer
-- coming soon ...
